netcdf 0103061300 {
dimensions:
	Num_Pireps = UNLIMITED ;
	Str1_Lngth = 9 ;
	Str2_Lngth = 8 ;
	Str3_Lngth = 1 ;
	Str4_Lngth = 256 ;
variables:
	int date(Num_Pireps) ;
		date:long_name = "Year/Month/Day of PIREP" ;
		date:units = "YYYYMMDD" ;
	short time(Num_Pireps) ;
		time:long_name = "Hour/Minute of PIREP" ;
		time:units = "HHMM" ;
	char rep_type(Num_Pireps, Str3_Lngth) ;
		rep_type:long_name = "Report Type" ;
		rep_type:units = "none" ;
		rep_type:valueP = "PIREP" ;
		rep_type:valueA = "AIREP" ;
	char acft(Num_Pireps, Str2_Lngth) ;
		acft:long_name = "Aircraft Type" ;
		acft:units = "none" ;
	float lat(Num_Pireps) ;
		lat:long_name = "Latitude of PIREP Location" ;
		lat:units = "Degrees North" ;
		lat:_FillValue = -99.f ;
	float lon(Num_Pireps) ;
		lon:long_name = "Longitude of PIREP Location" ;
		lon:units = "Degrees East" ;
		lon:_FillValue = -999.f ;
	int fl_level(Num_Pireps) ;
		fl_level:long_name = "Aircraft Flight Level" ;
		fl_level:units = "feet" ;
		fl_level:valid_range = 0, 60000 ;
		fl_level:_FillValue = -9 ;
	char pirep_type(Num_Pireps, Str3_Lngth) ;
		pirep_type:long_name = "PIREP Data Type" ;
		pirep_type:units = "none" ;
		pirep_type:valueN = "valid pirep with no mention of icing or turbulence." ;
		pirep_type:valueI = "icing data only (also clear above)." ;
		pirep_type:valueT = "turbulence data only." ;
		pirep_type:valueB = "both icing and turbulence data" ;
		pirep_type:valueC = "no icing or turbulence data, but clear skies" ;
		pirep_type:_FillValue = "N" ;
	int sky1_base(Num_Pireps) ;
		sky1_base:long_name = "Cloud Base" ;
		sky1_base:units = "feet" ;
		sky1_base:valid_range = 0, 60000 ;
		sky1_base:_FillValue = -9 ;
	int sky1_top(Num_Pireps) ;
		sky1_top:long_name = "Cloud Top" ;
		sky1_top:units = "feet" ;
		sky1_top:valid_range = 0, 60000 ;
		sky1_top:_FillValue = -9 ;
	short sky1_cg(Num_Pireps) ;
		sky1_cg:long_name = "Sky Coverage" ;
		sky1_cg:units = "none" ;
		sky1_cg:value-9 = "Not reported" ;
		sky1_cg:value0 = "CLEAR" ;
		sky1_cg:value1 = "-SCT" ;
		sky1_cg:value2 = "SCT" ;
		sky1_cg:value3 = "SCT-BKN" ;
		sky1_cg:value4 = "-BKN" ;
		sky1_cg:value5 = "BKN" ;
		sky1_cg:value6 = "BKN-OVC" ;
		sky1_cg:value7 = "-OVC" ;
		sky1_cg:value8 = "OVC" ;
		sky1_cg:value9 = "OBSCURD or WOXOF" ;
		sky1_cg:_FillValue = -9s ;
		sky1_cg:valid_range = 0s, 9s ;
	int sky2_base(Num_Pireps) ;
		sky2_base:long_name = "Cloud Base" ;
		sky2_base:units = "feet" ;
		sky2_base:valid_range = 0, 60000 ;
		sky2_base:_FillValue = -9 ;
	int sky2_top(Num_Pireps) ;
		sky2_top:long_name = "Cloud Top" ;
		sky2_top:units = "feet" ;
		sky2_top:valid_range = 0, 60000 ;
		sky2_top:_FillValue = -9 ;
	short sky2_cg(Num_Pireps) ;
		sky2_cg:long_name = "Sky Coverage" ;
		sky2_cg:units = "none" ;
		sky2_cg:value-9 = "Not reported" ;
		sky2_cg:value0 = "CLEAR" ;
		sky2_cg:value1 = "-SCT" ;
		sky2_cg:value2 = "SCT" ;
		sky2_cg:value3 = "SCT-BKN" ;
		sky2_cg:value4 = "-BKN" ;
		sky2_cg:value5 = "BKN" ;
		sky2_cg:value6 = "BKN-OVC" ;
		sky2_cg:value7 = "-OVC" ;
		sky2_cg:value8 = "OVC" ;
		sky2_cg:value9 = "OBSCURD or WOXOF" ;
		sky2_cg:_FillValue = -9s ;
		sky2_cg:valid_range = 0s, 9s ;
	int clr_abv(Num_Pireps) ;
		clr_abv:long_name = "Clear Above Level" ;
		clr_abv:units = "feet" ;
		clr_abv:valid_range = 0, 60000 ;
		clr_abv:_FillValue = -9 ;
	short wx_vs(Num_Pireps) ;
		wx_vs:long_name = "Visibility" ;
		wx_vs:units = "nautical miles" ;
		wx_vs:valid_range = 0s, 99s ;
		wx_vs:_FillValue = -9s ;
	short wx_ob(Num_Pireps) ;
		wx_ob:long_name = "Obstructions to Visibility" ;
		wx_ob:units = "none" ;
		wx_ob:value-9 = "Not reported" ;
		wx_ob:value2 = "VFR/GOOD/UNLIMITED" ;
		wx_ob:value3 = "CLEAR" ;
		wx_ob:value4 = "SMOKE" ;
		wx_ob:value5 = "HAZE" ;
		wx_ob:value6 = "DUST/ASH" ;
		wx_ob:value8 = "TORNADO" ;
		wx_ob:value9 = "SAND" ;
		wx_ob:value14 = "VIRGA" ;
		wx_ob:value17 = "LIGHTNING/THUNDERSTORM" ;
		wx_ob:value19 = "FUNNEL" ;
		wx_ob:value40 = "IFR/OBSCURED" ;
		wx_ob:value45 = "FOG/GROUND FOG" ;
		wx_ob:value48 = "FREEZING FOG" ;
		wx_ob:value51 = "DRIZZLE" ;
		wx_ob:value57 = "FREEZING DRIZZLE" ;
		wx_ob:value63 = "RAIN" ;
		wx_ob:value67 = "FREEZING RAIN" ;
		wx_ob:value73 = "SNOW" ;
		wx_ob:value77 = "GRAUPEL" ;
		wx_ob:value81 = "RAIN SHOWER" ;
		wx_ob:value86 = "SNOW SHOWER" ;
		wx_ob:value87 = "HAIL" ;
		wx_ob:valid_range = 0s, 99s ;
		wx_ob:_FillValue = -9s ;
	int wx_tmp(Num_Pireps) ;
		wx_tmp:long_name = "Temperature" ;
		wx_tmp:units = "degrees C" ;
		wx_tmp:valid_range = -200, 200 ;
		wx_tmp:_FillValue = -999 ;
	int wx_wdr(Num_Pireps) ;
		wx_wdr:long_name = "Wind Direction" ;
		wx_wdr:units = "degrees" ;
		wx_wdr:valid_range = 0, 359 ;
		wx_wdr:_FillValue = -9 ;
	int wx_wsp(Num_Pireps) ;
		wx_wsp:long_name = "Wind Speed" ;
		wx_wsp:units = "knots" ;
		wx_wsp:valid_range = 0, 999 ;
		wx_wsp:_FillValue = -9 ;
	int icg1_base(Num_Pireps) ;
		icg1_base:long_name = "Icing Base Flight Level" ;
		icg1_base:units = "feet" ;
		icg1_base:valid_range = 0, 60000 ;
		icg1_base:_FillValue = -9 ;
	int icg1_top(Num_Pireps) ;
		icg1_top:long_name = "Icing Top Flight Level" ;
		icg1_top:units = "feet" ;
		icg1_top:valid_range = 0, 60000 ;
		icg1_top:_FillValue = -9 ;
	short icg1_int(Num_Pireps) ;
		icg1_int:long_name = "Icing Intensity" ;
		icg1_int:units = "none" ;
		icg1_int:value-1 = "None" ;
		icg1_int:value1 = "Trace" ;
		icg1_int:value2 = "Trace to Light" ;
		icg1_int:value3 = "Light" ;
		icg1_int:value4 = "Light to Moderate" ;
		icg1_int:value5 = "Moderate" ;
		icg1_int:value6 = "Moderate to Heavy" ;
		icg1_int:value7 = "Heavy" ;
		icg1_int:value8 = "Severe" ;
		icg1_int:_FillValue = -9s ;
	short icg1_type(Num_Pireps) ;
		icg1_type:long_name = "Icing Type" ;
		icg1_type:units = "none" ;
		icg1_type:value1 = "Rime" ;
		icg1_type:value2 = "Clear" ;
		icg1_type:value3 = "Mixed" ;
		icg1_type:_FillValue = -9s ;
	int icg2_base(Num_Pireps) ;
		icg2_base:long_name = "Icing Base Flight Level" ;
		icg2_base:units = "feet" ;
		icg2_base:valid_range = 0, 60000 ;
		icg2_base:_FillValue = -9 ;
	int icg2_top(Num_Pireps) ;
		icg2_top:long_name = "Icing Top Flight Level" ;
		icg2_top:units = "feet" ;
		icg2_top:valid_range = 0, 60000 ;
		icg2_top:_FillValue = -9 ;
	short icg2_int(Num_Pireps) ;
		icg2_int:long_name = "Icing Intensity" ;
		icg2_int:units = "none" ;
		icg2_int:value-1 = "None" ;
		icg2_int:value1 = "Trace" ;
		icg2_int:value2 = "Trace to Light" ;
		icg2_int:value3 = "Light" ;
		icg2_int:value4 = "Light to Moderate" ;
		icg2_int:value5 = "Moderate" ;
		icg2_int:value6 = "Moderate to Heavy" ;
		icg2_int:value7 = "Heavy" ;
		icg2_int:value8 = "Severe" ;
		icg2_int:_FillValue = -9s ;
	short icg2_type(Num_Pireps) ;
		icg2_type:long_name = "Icing Type" ;
		icg2_type:units = "none" ;
		icg2_type:value1 = "Rime" ;
		icg2_type:value2 = "Clear" ;
		icg2_type:value3 = "Mixed" ;
		icg2_type:_FillValue = -9s ;
	int trb1_base(Num_Pireps) ;
		trb1_base:long_name = "Turbulence Base Flight Level" ;
		trb1_base:units = "feet" ;
		trb1_base:valid_range = 0, 60000 ;
		trb1_base:_FillValue = -9 ;
	int trb1_top(Num_Pireps) ;
		trb1_top:long_name = "Turbulence Top Flight Level" ;
		trb1_top:units = "feet" ;
		trb1_top:valid_range = 0, 60000 ;
		trb1_top:_FillValue = -9 ;
	short trb1_frq(Num_Pireps) ;
		trb1_frq:long_name = "Turbulence Frequency" ;
		trb1_frq:units = "none" ;
		trb1_frq:value1 = "Occasional" ;
		trb1_frq:value2 = "Intermittent" ;
		trb1_frq:value3 = "Continuous" ;
		trb1_frq:_FillValue = -9s ;
	short trb1_int(Num_Pireps) ;
		trb1_int:long_name = "Turbulence Intensity" ;
		trb1_int:units = "none" ;
		trb1_int:value0 = "None/Smooth" ;
		trb1_int:value1 = "Smooth to Light" ;
		trb1_int:value2 = "Light to Moderate" ;
		trb1_int:value3 = "Moderate" ;
		trb1_int:value4 = "Moderate to Severe" ;
		trb1_int:value5 = "Severe" ;
		trb1_int:value6 = "Severe to Extreme" ;
		trb1_int:value7 = "Extreme" ;
		trb1_int:_FillValue = -9s ;
	short trb1_type(Num_Pireps) ;
		trb1_type:long_name = "Turbulence Type" ;
		trb1_type:units = "none" ;
		trb1_type:value1 = "Chop" ;
		trb1_type:value2 = "Clear Air Turbulence" ;
		trb1_type:value3 = "Low-level Wind Shear" ;
		trb1_type:value4 = "MTN Wave" ;
		trb1_type:_FillValue = -9s ;
	int trb2_base(Num_Pireps) ;
		trb2_base:long_name = "Turbulence Base Flight Level" ;
		trb2_base:units = "feet" ;
		trb2_base:valid_range = 0, 60000 ;
		trb2_base:_FillValue = -9 ;
	int trb2_top(Num_Pireps) ;
		trb2_top:long_name = "Turbulence Top Flight Level" ;
		trb2_top:units = "feet" ;
		trb2_top:valid_range = 0, 60000 ;
		trb2_top:_FillValue = -9 ;
	short trb2_frq(Num_Pireps) ;
		trb2_frq:long_name = "Turbulence Frequency" ;
		trb2_frq:units = "none" ;
		trb2_frq:value1 = "Occasional" ;
		trb2_frq:value2 = "Intermittent" ;
		trb2_frq:value3 = "Continuous" ;
		trb2_frq:_FillValue = -9s ;
	short trb2_int(Num_Pireps) ;
		trb2_int:long_name = "Turbulence Intensity" ;
		trb2_int:units = "none" ;
		trb2_int:value0 = "None/Smooth" ;
		trb2_int:value1 = "Smooth to Light" ;
		trb2_int:value2 = "Light to Moderate" ;
		trb2_int:value3 = "Moderate" ;
		trb2_int:value4 = "Moderate to Severe" ;
		trb2_int:value5 = "Severe" ;
		trb2_int:value6 = "Severe to Extreme" ;
		trb2_int:value7 = "Extreme" ;
		trb2_int:_FillValue = -9s ;
	short trb2_type(Num_Pireps) ;
		trb2_type:long_name = "Turbulence Type" ;
		trb2_type:units = "none" ;
		trb2_type:value1 = "Chop" ;
		trb2_type:value2 = "Clear Air Turbulence" ;
		trb2_type:value3 = "Low-level Wind Shear" ;
		trb2_type:value4 = "MTN Wave" ;
		trb2_type:_FillValue = -9s ;
	char raw_pirep(Num_Pireps, Str4_Lngth) ;
		raw_pirep:long_name = "Raw Pirep" ;

// global attributes:
		:Title = "Decoded PIREPs/AIREPs" ;
                :Version = "2.2a";
}
